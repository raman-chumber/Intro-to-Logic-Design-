module orgate(in1, in2, out);
input in1, in2;
output out;

wire in1, in2, out;

or g1(out, in1, in2, out);

endmodule